-- DE0_CV_QSYS.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DE0_CV_QSYS is
	port (
		clk_clk                 : in    std_logic                     := '0';             --              clk.clk
		clk_sdram_clk           : out   std_logic;                                        --        clk_sdram.clk
		keys_wire_export        : in    std_logic_vector(3 downto 0)  := (others => '0'); --        keys_wire.export
		leds_wire_export        : out   std_logic_vector(9 downto 0);                     --        leds_wire.export
		line_export             : out   std_logic;                                        --             line.export
		pll_locked_export       : out   std_logic;                                        --       pll_locked.export
		reset_reset_n           : in    std_logic                     := '0';             --            reset.reset_n
		sdram_wire_addr         : out   std_logic_vector(12 downto 0);                    --       sdram_wire.addr
		sdram_wire_ba           : out   std_logic_vector(1 downto 0);                     --                 .ba
		sdram_wire_cas_n        : out   std_logic;                                        --                 .cas_n
		sdram_wire_cke          : out   std_logic;                                        --                 .cke
		sdram_wire_cs_n         : out   std_logic;                                        --                 .cs_n
		sdram_wire_dq           : inout std_logic_vector(15 downto 0) := (others => '0'); --                 .dq
		sdram_wire_dqm          : out   std_logic_vector(1 downto 0);                     --                 .dqm
		sdram_wire_ras_n        : out   std_logic;                                        --                 .ras_n
		sdram_wire_we_n         : out   std_logic;                                        --                 .we_n
		seg7_digits_wire_export : out   std_logic_vector(23 downto 0);                    -- seg7_digits_wire.export
		switches_wire_export    : in    std_logic_vector(9 downto 0)  := (others => '0')  --    switches_wire.export
	);
end entity DE0_CV_QSYS;

architecture rtl of DE0_CV_QSYS is
	component DE0_CV_QSYS_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component DE0_CV_QSYS_jtag_uart;

	component DE0_CV_QSYS_keys is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component DE0_CV_QSYS_keys;

	component DE0_CV_QSYS_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component DE0_CV_QSYS_leds;

	component altera_avalon_mm_clock_crossing_bridge is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			HDL_ADDR_WIDTH      : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             -- clk
			m0_reset         : in  std_logic                     := 'X';             -- reset
			s0_clk           : in  std_logic                     := 'X';             -- clk
			s0_reset         : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(11 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component altera_avalon_mm_clock_crossing_bridge;

	component DE0_CV_QSYS_nios2_qsys is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component DE0_CV_QSYS_nios2_qsys;

	component DE0_CV_QSYS_onchip_mem is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component DE0_CV_QSYS_onchip_mem;

	component DE0_CV_QSYS_pll is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component DE0_CV_QSYS_pll;

	component DE0_CV_QSYS_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component DE0_CV_QSYS_sdram;

	component DE0_CV_QSYS_seg7_digits is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(23 downto 0)                     -- export
		);
	end component DE0_CV_QSYS_seg7_digits;

	component DE0_CV_QSYS_switches is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component DE0_CV_QSYS_switches;

	component DE0_CV_QSYS_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component DE0_CV_QSYS_sysid_qsys;

	component DE0_CV_QSYS_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component DE0_CV_QSYS_timer;

	component eln is
		port (
			rd        : in  std_logic                    := 'X';             -- read
			wr        : in  std_logic                    := 'X';             -- write
			D_in      : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			D_out     : out std_logic_vector(7 downto 0);                    -- readdata
			Addr      : in  std_logic_vector(1 downto 0) := (others => 'X'); -- address
			Clk       : in  std_logic                    := 'X';             -- clk
			reset_n   : in  std_logic                    := 'X';             -- reset_n
			IRQ_ELN_n : out std_logic;                                       -- irq_n
			Line_ELN  : out std_logic                                        -- export
		);
	end component eln;

	component DE0_CV_QSYS_mm_interconnect_0 is
		port (
			pll_outclk0_clk                              : in  std_logic                     := 'X';             -- clk
			nios2_qsys_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_qsys_data_master_address               : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_qsys_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2_qsys_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_qsys_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios2_qsys_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_data_master_readdatavalid         : out std_logic;                                        -- readdatavalid
			nios2_qsys_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios2_qsys_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_qsys_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios2_qsys_instruction_master_address        : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_qsys_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios2_qsys_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios2_qsys_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_instruction_master_readdatavalid  : out std_logic;                                        -- readdatavalid
			jtag_uart_avalon_jtag_slave_address          : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write            : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read             : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect       : out std_logic;                                        -- chipselect
			mm_clock_crossing_bridge_0_s0_address        : out std_logic_vector(11 downto 0);                    -- address
			mm_clock_crossing_bridge_0_s0_write          : out std_logic;                                        -- write
			mm_clock_crossing_bridge_0_s0_read           : out std_logic;                                        -- read
			mm_clock_crossing_bridge_0_s0_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mm_clock_crossing_bridge_0_s0_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			mm_clock_crossing_bridge_0_s0_burstcount     : out std_logic_vector(0 downto 0);                     -- burstcount
			mm_clock_crossing_bridge_0_s0_byteenable     : out std_logic_vector(3 downto 0);                     -- byteenable
			mm_clock_crossing_bridge_0_s0_readdatavalid  : in  std_logic                     := 'X';             -- readdatavalid
			mm_clock_crossing_bridge_0_s0_waitrequest    : in  std_logic                     := 'X';             -- waitrequest
			mm_clock_crossing_bridge_0_s0_debugaccess    : out std_logic;                                        -- debugaccess
			nios2_qsys_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_qsys_debug_mem_slave_write             : out std_logic;                                        -- write
			nios2_qsys_debug_mem_slave_read              : out std_logic;                                        -- read
			nios2_qsys_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_qsys_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_qsys_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_qsys_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_qsys_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			onchip_mem_s1_address                        : out std_logic_vector(14 downto 0);                    -- address
			onchip_mem_s1_write                          : out std_logic;                                        -- write
			onchip_mem_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_mem_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_mem_s1_byteenable                     : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_mem_s1_chipselect                     : out std_logic;                                        -- chipselect
			onchip_mem_s1_clken                          : out std_logic;                                        -- clken
			sdram_s1_address                             : out std_logic_vector(24 downto 0);                    -- address
			sdram_s1_write                               : out std_logic;                                        -- write
			sdram_s1_read                                : out std_logic;                                        -- read
			sdram_s1_readdata                            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                           : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                          : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                          : out std_logic                                         -- chipselect
		);
	end component DE0_CV_QSYS_mm_interconnect_0;

	component DE0_CV_QSYS_mm_interconnect_1 is
		port (
			pll_outclk2_clk                                                 : in  std_logic                     := 'X';             -- clk
			mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			transmitter_reset_n_reset_bridge_in_reset_reset                 : in  std_logic                     := 'X';             -- reset
			mm_clock_crossing_bridge_0_m0_address                           : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			mm_clock_crossing_bridge_0_m0_waitrequest                       : out std_logic;                                        -- waitrequest
			mm_clock_crossing_bridge_0_m0_burstcount                        : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			mm_clock_crossing_bridge_0_m0_byteenable                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			mm_clock_crossing_bridge_0_m0_read                              : in  std_logic                     := 'X';             -- read
			mm_clock_crossing_bridge_0_m0_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			mm_clock_crossing_bridge_0_m0_readdatavalid                     : out std_logic;                                        -- readdatavalid
			mm_clock_crossing_bridge_0_m0_write                             : in  std_logic                     := 'X';             -- write
			mm_clock_crossing_bridge_0_m0_writedata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			mm_clock_crossing_bridge_0_m0_debugaccess                       : in  std_logic                     := 'X';             -- debugaccess
			keys_s1_address                                                 : out std_logic_vector(1 downto 0);                     -- address
			keys_s1_write                                                   : out std_logic;                                        -- write
			keys_s1_readdata                                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			keys_s1_writedata                                               : out std_logic_vector(31 downto 0);                    -- writedata
			keys_s1_chipselect                                              : out std_logic;                                        -- chipselect
			leds_s1_address                                                 : out std_logic_vector(2 downto 0);                     -- address
			leds_s1_write                                                   : out std_logic;                                        -- write
			leds_s1_readdata                                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_s1_writedata                                               : out std_logic_vector(31 downto 0);                    -- writedata
			leds_s1_chipselect                                              : out std_logic;                                        -- chipselect
			seg7_digits_s1_address                                          : out std_logic_vector(2 downto 0);                     -- address
			seg7_digits_s1_write                                            : out std_logic;                                        -- write
			seg7_digits_s1_readdata                                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			seg7_digits_s1_writedata                                        : out std_logic_vector(31 downto 0);                    -- writedata
			seg7_digits_s1_chipselect                                       : out std_logic;                                        -- chipselect
			switches_s1_address                                             : out std_logic_vector(1 downto 0);                     -- address
			switches_s1_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sysid_qsys_control_slave_address                                : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_control_slave_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_s1_address                                                : out std_logic_vector(2 downto 0);                     -- address
			timer_s1_write                                                  : out std_logic;                                        -- write
			timer_s1_readdata                                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_s1_writedata                                              : out std_logic_vector(15 downto 0);                    -- writedata
			timer_s1_chipselect                                             : out std_logic;                                        -- chipselect
			transmitter_avalon_eln_address                                  : out std_logic_vector(1 downto 0);                     -- address
			transmitter_avalon_eln_write                                    : out std_logic;                                        -- write
			transmitter_avalon_eln_read                                     : out std_logic;                                        -- read
			transmitter_avalon_eln_readdata                                 : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			transmitter_avalon_eln_writedata                                : out std_logic_vector(7 downto 0)                      -- writedata
		);
	end component DE0_CV_QSYS_mm_interconnect_1;

	component DE0_CV_QSYS_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component DE0_CV_QSYS_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component de0_cv_qsys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component de0_cv_qsys_rst_controller;

	component de0_cv_qsys_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component de0_cv_qsys_rst_controller_001;

	signal pll_outclk0_clk                                               : std_logic;                     -- pll:outclk_0 -> [irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, jtag_uart:clk, mm_clock_crossing_bridge_0:s0_clk, mm_interconnect_0:pll_outclk0_clk, nios2_qsys:clk, onchip_mem:clk, rst_controller:clk, sdram:clk]
	signal pll_outclk2_clk                                               : std_logic;                     -- pll:outclk_2 -> [irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, keys:clk, leds:clk, mm_clock_crossing_bridge_0:m0_clk, mm_interconnect_1:pll_outclk2_clk, rst_controller_001:clk, seg7_digits:clk, switches:clk, sysid_qsys:clock, timer:clk, transmitter:Clk]
	signal nios2_qsys_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	signal nios2_qsys_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	signal nios2_qsys_data_master_debugaccess                            : std_logic;                     -- nios2_qsys:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	signal nios2_qsys_data_master_address                                : std_logic_vector(26 downto 0); -- nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	signal nios2_qsys_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	signal nios2_qsys_data_master_read                                   : std_logic;                     -- nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	signal nios2_qsys_data_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:nios2_qsys_data_master_readdatavalid -> nios2_qsys:d_readdatavalid
	signal nios2_qsys_data_master_write                                  : std_logic;                     -- nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	signal nios2_qsys_data_master_writedata                              : std_logic_vector(31 downto 0); -- nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	signal nios2_qsys_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	signal nios2_qsys_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	signal nios2_qsys_instruction_master_address                         : std_logic_vector(26 downto 0); -- nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	signal nios2_qsys_instruction_master_read                            : std_logic;                     -- nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	signal nios2_qsys_instruction_master_readdatavalid                   : std_logic;                     -- mm_interconnect_0:nios2_qsys_instruction_master_readdatavalid -> nios2_qsys:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata         : std_logic_vector(31 downto 0); -- nios2_qsys:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest      : std_logic;                     -- nios2_qsys:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess      : std_logic;                     -- mm_interconnect_0:nios2_qsys_debug_mem_slave_debugaccess -> nios2_qsys:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_qsys_debug_mem_slave_address -> nios2_qsys:debug_mem_slave_address
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_read             : std_logic;                     -- mm_interconnect_0:nios2_qsys_debug_mem_slave_read -> nios2_qsys:debug_mem_slave_read
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_qsys_debug_mem_slave_byteenable -> nios2_qsys:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_write            : std_logic;                     -- mm_interconnect_0:nios2_qsys_debug_mem_slave_write -> nios2_qsys:debug_mem_slave_write
	signal mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_debug_mem_slave_writedata -> nios2_qsys:debug_mem_slave_writedata
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata      : std_logic_vector(31 downto 0); -- mm_clock_crossing_bridge_0:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdata
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest   : std_logic;                     -- mm_clock_crossing_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_waitrequest
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess   : std_logic;                     -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_debugaccess -> mm_clock_crossing_bridge_0:s0_debugaccess
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address       : std_logic_vector(11 downto 0); -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_address -> mm_clock_crossing_bridge_0:s0_address
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read          : std_logic;                     -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_read -> mm_clock_crossing_bridge_0:s0_read
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_byteenable -> mm_clock_crossing_bridge_0:s0_byteenable
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid : std_logic;                     -- mm_clock_crossing_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdatavalid
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write         : std_logic;                     -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_write -> mm_clock_crossing_bridge_0:s0_write
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_writedata -> mm_clock_crossing_bridge_0:s0_writedata
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_burstcount -> mm_clock_crossing_bridge_0:s0_burstcount
	signal mm_interconnect_0_onchip_mem_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_chipselect -> onchip_mem:chipselect
	signal mm_interconnect_0_onchip_mem_s1_readdata                      : std_logic_vector(31 downto 0); -- onchip_mem:readdata -> mm_interconnect_0:onchip_mem_s1_readdata
	signal mm_interconnect_0_onchip_mem_s1_address                       : std_logic_vector(14 downto 0); -- mm_interconnect_0:onchip_mem_s1_address -> onchip_mem:address
	signal mm_interconnect_0_onchip_mem_s1_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_mem_s1_byteenable -> onchip_mem:byteenable
	signal mm_interconnect_0_onchip_mem_s1_write                         : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_write -> onchip_mem:write
	signal mm_interconnect_0_onchip_mem_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_mem_s1_writedata -> onchip_mem:writedata
	signal mm_interconnect_0_onchip_mem_s1_clken                         : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_clken -> onchip_mem:clken
	signal mm_interconnect_0_sdram_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                           : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                        : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                            : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                               : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                      : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                              : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_clock_crossing_bridge_0_m0_waitrequest                     : std_logic;                     -- mm_interconnect_1:mm_clock_crossing_bridge_0_m0_waitrequest -> mm_clock_crossing_bridge_0:m0_waitrequest
	signal mm_clock_crossing_bridge_0_m0_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_1:mm_clock_crossing_bridge_0_m0_readdata -> mm_clock_crossing_bridge_0:m0_readdata
	signal mm_clock_crossing_bridge_0_m0_debugaccess                     : std_logic;                     -- mm_clock_crossing_bridge_0:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_debugaccess
	signal mm_clock_crossing_bridge_0_m0_address                         : std_logic_vector(11 downto 0); -- mm_clock_crossing_bridge_0:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_address
	signal mm_clock_crossing_bridge_0_m0_read                            : std_logic;                     -- mm_clock_crossing_bridge_0:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_read
	signal mm_clock_crossing_bridge_0_m0_byteenable                      : std_logic_vector(3 downto 0);  -- mm_clock_crossing_bridge_0:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_byteenable
	signal mm_clock_crossing_bridge_0_m0_readdatavalid                   : std_logic;                     -- mm_interconnect_1:mm_clock_crossing_bridge_0_m0_readdatavalid -> mm_clock_crossing_bridge_0:m0_readdatavalid
	signal mm_clock_crossing_bridge_0_m0_writedata                       : std_logic_vector(31 downto 0); -- mm_clock_crossing_bridge_0:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_writedata
	signal mm_clock_crossing_bridge_0_m0_write                           : std_logic;                     -- mm_clock_crossing_bridge_0:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_write
	signal mm_clock_crossing_bridge_0_m0_burstcount                      : std_logic_vector(0 downto 0);  -- mm_clock_crossing_bridge_0:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_burstcount
	signal mm_interconnect_1_transmitter_avalon_eln_readdata             : std_logic_vector(7 downto 0);  -- transmitter:D_out -> mm_interconnect_1:transmitter_avalon_eln_readdata
	signal mm_interconnect_1_transmitter_avalon_eln_address              : std_logic_vector(1 downto 0);  -- mm_interconnect_1:transmitter_avalon_eln_address -> transmitter:Addr
	signal mm_interconnect_1_transmitter_avalon_eln_read                 : std_logic;                     -- mm_interconnect_1:transmitter_avalon_eln_read -> transmitter:rd
	signal mm_interconnect_1_transmitter_avalon_eln_write                : std_logic;                     -- mm_interconnect_1:transmitter_avalon_eln_write -> transmitter:wr
	signal mm_interconnect_1_transmitter_avalon_eln_writedata            : std_logic_vector(7 downto 0);  -- mm_interconnect_1:transmitter_avalon_eln_writedata -> transmitter:D_in
	signal mm_interconnect_1_sysid_qsys_control_slave_readdata           : std_logic_vector(31 downto 0); -- sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	signal mm_interconnect_1_sysid_qsys_control_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	signal mm_interconnect_1_timer_s1_chipselect                         : std_logic;                     -- mm_interconnect_1:timer_s1_chipselect -> timer:chipselect
	signal mm_interconnect_1_timer_s1_readdata                           : std_logic_vector(15 downto 0); -- timer:readdata -> mm_interconnect_1:timer_s1_readdata
	signal mm_interconnect_1_timer_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_1:timer_s1_address -> timer:address
	signal mm_interconnect_1_timer_s1_write                              : std_logic;                     -- mm_interconnect_1:timer_s1_write -> mm_interconnect_1_timer_s1_write:in
	signal mm_interconnect_1_timer_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_1:timer_s1_writedata -> timer:writedata
	signal mm_interconnect_1_keys_s1_chipselect                          : std_logic;                     -- mm_interconnect_1:keys_s1_chipselect -> keys:chipselect
	signal mm_interconnect_1_keys_s1_readdata                            : std_logic_vector(31 downto 0); -- keys:readdata -> mm_interconnect_1:keys_s1_readdata
	signal mm_interconnect_1_keys_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_1:keys_s1_address -> keys:address
	signal mm_interconnect_1_keys_s1_write                               : std_logic;                     -- mm_interconnect_1:keys_s1_write -> mm_interconnect_1_keys_s1_write:in
	signal mm_interconnect_1_keys_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_1:keys_s1_writedata -> keys:writedata
	signal mm_interconnect_1_switches_s1_readdata                        : std_logic_vector(31 downto 0); -- switches:readdata -> mm_interconnect_1:switches_s1_readdata
	signal mm_interconnect_1_switches_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_1:switches_s1_address -> switches:address
	signal mm_interconnect_1_leds_s1_chipselect                          : std_logic;                     -- mm_interconnect_1:leds_s1_chipselect -> leds:chipselect
	signal mm_interconnect_1_leds_s1_readdata                            : std_logic_vector(31 downto 0); -- leds:readdata -> mm_interconnect_1:leds_s1_readdata
	signal mm_interconnect_1_leds_s1_address                             : std_logic_vector(2 downto 0);  -- mm_interconnect_1:leds_s1_address -> leds:address
	signal mm_interconnect_1_leds_s1_write                               : std_logic;                     -- mm_interconnect_1:leds_s1_write -> mm_interconnect_1_leds_s1_write:in
	signal mm_interconnect_1_leds_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_1:leds_s1_writedata -> leds:writedata
	signal mm_interconnect_1_seg7_digits_s1_chipselect                   : std_logic;                     -- mm_interconnect_1:seg7_digits_s1_chipselect -> seg7_digits:chipselect
	signal mm_interconnect_1_seg7_digits_s1_readdata                     : std_logic_vector(31 downto 0); -- seg7_digits:readdata -> mm_interconnect_1:seg7_digits_s1_readdata
	signal mm_interconnect_1_seg7_digits_s1_address                      : std_logic_vector(2 downto 0);  -- mm_interconnect_1:seg7_digits_s1_address -> seg7_digits:address
	signal mm_interconnect_1_seg7_digits_s1_write                        : std_logic;                     -- mm_interconnect_1:seg7_digits_s1_write -> mm_interconnect_1_seg7_digits_s1_write:in
	signal mm_interconnect_1_seg7_digits_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_1:seg7_digits_s1_writedata -> seg7_digits:writedata
	signal irq_mapper_receiver2_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver2_irq
	signal nios2_qsys_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_qsys:irq
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal transmitter_irq_eln_n_irq                                     : std_logic;                     -- transmitter:IRQ_ELN_n -> transmitter_irq_eln_n_irq:in
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	signal irq_synchronizer_001_receiver_irq                             : std_logic_vector(0 downto 0);  -- timer:irq -> irq_synchronizer_001:receiver_irq
	signal irq_mapper_receiver3_irq                                      : std_logic;                     -- irq_synchronizer_002:sender_irq -> irq_mapper:receiver3_irq
	signal irq_synchronizer_002_receiver_irq                             : std_logic_vector(0 downto 0);  -- keys:irq -> irq_synchronizer_002:receiver_irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, mm_clock_crossing_bridge_0:s0_reset, mm_interconnect_0:nios2_qsys_reset_reset_bridge_in_reset_reset, onchip_mem:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [nios2_qsys:reset_req, onchip_mem:reset_req, rst_translator:reset_req_in]
	signal nios2_qsys_debug_reset_request_reset                          : std_logic;                     -- nios2_qsys:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, mm_clock_crossing_bridge_0:m0_reset, mm_interconnect_1:mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:transmitter_reset_n_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset                            : std_logic;                     -- rst_controller_002:reset_out -> rst_controller_002_reset_out_reset:in
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [pll:rst, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                     : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv               : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_1_timer_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_1_timer_s1_write:inv -> timer:write_n
	signal mm_interconnect_1_keys_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_1_keys_s1_write:inv -> keys:write_n
	signal mm_interconnect_1_leds_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_1_leds_s1_write:inv -> leds:write_n
	signal mm_interconnect_1_seg7_digits_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_1_seg7_digits_s1_write:inv -> seg7_digits:write_n
	signal irq_synchronizer_receiver_inv                                 : std_logic_vector(0 downto 0);  -- transmitter_irq_eln_n_irq:inv -> irq_synchronizer:receiver_irq
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [jtag_uart:rst_n, nios2_qsys:reset_n, sdram:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [keys:reset_n, leds:reset_n, seg7_digits:reset_n, switches:reset_n, sysid_qsys:reset_n, timer:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> transmitter:reset_n

begin

	jtag_uart : component DE0_CV_QSYS_jtag_uart
		port map (
			clk            => pll_outclk0_clk,                                               --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver2_irq                                       --               irq.irq
		);

	keys : component DE0_CV_QSYS_keys
		port map (
			clk        => pll_outclk2_clk,                              --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_keys_s1_address,            --                  s1.address
			write_n    => mm_interconnect_1_keys_s1_write_ports_inv,    --                    .write_n
			writedata  => mm_interconnect_1_keys_s1_writedata,          --                    .writedata
			chipselect => mm_interconnect_1_keys_s1_chipselect,         --                    .chipselect
			readdata   => mm_interconnect_1_keys_s1_readdata,           --                    .readdata
			in_port    => keys_wire_export,                             -- external_connection.export
			irq        => irq_synchronizer_002_receiver_irq(0)          --                 irq.irq
		);

	leds : component DE0_CV_QSYS_leds
		port map (
			clk        => pll_outclk2_clk,                              --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_leds_s1_address,            --                  s1.address
			write_n    => mm_interconnect_1_leds_s1_write_ports_inv,    --                    .write_n
			writedata  => mm_interconnect_1_leds_s1_writedata,          --                    .writedata
			chipselect => mm_interconnect_1_leds_s1_chipselect,         --                    .chipselect
			readdata   => mm_interconnect_1_leds_s1_readdata,           --                    .readdata
			out_port   => leds_wire_export                              -- external_connection.export
		);

	mm_clock_crossing_bridge_0 : component altera_avalon_mm_clock_crossing_bridge
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			HDL_ADDR_WIDTH      => 12,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 4,
			RESPONSE_FIFO_DEPTH => 4,
			MASTER_SYNC_DEPTH   => 2,
			SLAVE_SYNC_DEPTH    => 2
		)
		port map (
			m0_clk           => pll_outclk2_clk,                                               --   m0_clk.clk
			m0_reset         => rst_controller_001_reset_out_reset,                            -- m0_reset.reset
			s0_clk           => pll_outclk0_clk,                                               --   s0_clk.clk
			s0_reset         => rst_controller_reset_out_reset,                                -- s0_reset.reset
			s0_waitrequest   => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest,   --       s0.waitrequest
			s0_readdata      => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata,      --         .readdata
			s0_readdatavalid => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid, --         .readdatavalid
			s0_burstcount    => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount,    --         .burstcount
			s0_writedata     => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata,     --         .writedata
			s0_address       => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address,       --         .address
			s0_write         => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write,         --         .write
			s0_read          => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read,          --         .read
			s0_byteenable    => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable,    --         .byteenable
			s0_debugaccess   => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess,   --         .debugaccess
			m0_waitrequest   => mm_clock_crossing_bridge_0_m0_waitrequest,                     --       m0.waitrequest
			m0_readdata      => mm_clock_crossing_bridge_0_m0_readdata,                        --         .readdata
			m0_readdatavalid => mm_clock_crossing_bridge_0_m0_readdatavalid,                   --         .readdatavalid
			m0_burstcount    => mm_clock_crossing_bridge_0_m0_burstcount,                      --         .burstcount
			m0_writedata     => mm_clock_crossing_bridge_0_m0_writedata,                       --         .writedata
			m0_address       => mm_clock_crossing_bridge_0_m0_address,                         --         .address
			m0_write         => mm_clock_crossing_bridge_0_m0_write,                           --         .write
			m0_read          => mm_clock_crossing_bridge_0_m0_read,                            --         .read
			m0_byteenable    => mm_clock_crossing_bridge_0_m0_byteenable,                      --         .byteenable
			m0_debugaccess   => mm_clock_crossing_bridge_0_m0_debugaccess                      --         .debugaccess
		);

	nios2_qsys : component DE0_CV_QSYS_nios2_qsys
		port map (
			clk                                 => pll_outclk0_clk,                                          --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                 --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                       --                          .reset_req
			d_address                           => nios2_qsys_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_qsys_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_qsys_data_master_read,                              --                          .read
			d_readdata                          => nios2_qsys_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_qsys_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_qsys_data_master_write,                             --                          .write
			d_writedata                         => nios2_qsys_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_qsys_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_qsys_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_qsys_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_qsys_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_qsys_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_qsys_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_qsys_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_qsys_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_qsys_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_qsys_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_qsys_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_qsys_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                      -- custom_instruction_master.readra
		);

	onchip_mem : component DE0_CV_QSYS_onchip_mem
		port map (
			clk        => pll_outclk0_clk,                            --   clk1.clk
			address    => mm_interconnect_0_onchip_mem_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_mem_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_mem_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_mem_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_mem_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_mem_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_mem_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,         --       .reset_req
			freeze     => '0'                                         -- (terminated)
		);

	pll : component DE0_CV_QSYS_pll
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_outclk0_clk,         -- outclk0.clk
			outclk_1 => clk_sdram_clk,           -- outclk1.clk
			outclk_2 => pll_outclk2_clk,         -- outclk2.clk
			locked   => pll_locked_export        --  locked.export
		);

	sdram : component DE0_CV_QSYS_sdram
		port map (
			clk            => pll_outclk0_clk,                                 --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	seg7_digits : component DE0_CV_QSYS_seg7_digits
		port map (
			clk        => pll_outclk2_clk,                                  --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_1_seg7_digits_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_seg7_digits_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_seg7_digits_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_seg7_digits_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_seg7_digits_s1_readdata,        --                    .readdata
			out_port   => seg7_digits_wire_export                           -- external_connection.export
		);

	switches : component DE0_CV_QSYS_switches
		port map (
			clk      => pll_outclk2_clk,                              --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_1_switches_s1_address,        --                  s1.address
			readdata => mm_interconnect_1_switches_s1_readdata,       --                    .readdata
			in_port  => switches_wire_export                          -- external_connection.export
		);

	sysid_qsys : component DE0_CV_QSYS_sysid_qsys
		port map (
			clock    => pll_outclk2_clk,                                       --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,          --         reset.reset_n
			readdata => mm_interconnect_1_sysid_qsys_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_1_sysid_qsys_control_slave_address(0)  --              .address
		);

	timer : component DE0_CV_QSYS_timer
		port map (
			clk        => pll_outclk2_clk,                              --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_1_timer_s1_address,           --    s1.address
			writedata  => mm_interconnect_1_timer_s1_writedata,         --      .writedata
			readdata   => mm_interconnect_1_timer_s1_readdata,          --      .readdata
			chipselect => mm_interconnect_1_timer_s1_chipselect,        --      .chipselect
			write_n    => mm_interconnect_1_timer_s1_write_ports_inv,   --      .write_n
			irq        => irq_synchronizer_001_receiver_irq(0)          --   irq.irq
		);

	transmitter : component eln
		port map (
			rd        => mm_interconnect_1_transmitter_avalon_eln_read,      -- avalon_eln.read
			wr        => mm_interconnect_1_transmitter_avalon_eln_write,     --           .write
			D_in      => mm_interconnect_1_transmitter_avalon_eln_writedata, --           .writedata
			D_out     => mm_interconnect_1_transmitter_avalon_eln_readdata,  --           .readdata
			Addr      => mm_interconnect_1_transmitter_avalon_eln_address,   --           .address
			Clk       => pll_outclk2_clk,                                    --      clock.clk
			reset_n   => rst_controller_002_reset_out_reset_ports_inv,       --    reset_n.reset_n
			IRQ_ELN_n => transmitter_irq_eln_n_irq,                          --  Irq_ELN_n.irq_n
			Line_ELN  => line_export                                         --       Line.export
		);

	mm_interconnect_0 : component DE0_CV_QSYS_mm_interconnect_0
		port map (
			pll_outclk0_clk                              => pll_outclk0_clk,                                               --                            pll_outclk0.clk
			nios2_qsys_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                -- nios2_qsys_reset_reset_bridge_in_reset.reset
			nios2_qsys_data_master_address               => nios2_qsys_data_master_address,                                --                 nios2_qsys_data_master.address
			nios2_qsys_data_master_waitrequest           => nios2_qsys_data_master_waitrequest,                            --                                       .waitrequest
			nios2_qsys_data_master_byteenable            => nios2_qsys_data_master_byteenable,                             --                                       .byteenable
			nios2_qsys_data_master_read                  => nios2_qsys_data_master_read,                                   --                                       .read
			nios2_qsys_data_master_readdata              => nios2_qsys_data_master_readdata,                               --                                       .readdata
			nios2_qsys_data_master_readdatavalid         => nios2_qsys_data_master_readdatavalid,                          --                                       .readdatavalid
			nios2_qsys_data_master_write                 => nios2_qsys_data_master_write,                                  --                                       .write
			nios2_qsys_data_master_writedata             => nios2_qsys_data_master_writedata,                              --                                       .writedata
			nios2_qsys_data_master_debugaccess           => nios2_qsys_data_master_debugaccess,                            --                                       .debugaccess
			nios2_qsys_instruction_master_address        => nios2_qsys_instruction_master_address,                         --          nios2_qsys_instruction_master.address
			nios2_qsys_instruction_master_waitrequest    => nios2_qsys_instruction_master_waitrequest,                     --                                       .waitrequest
			nios2_qsys_instruction_master_read           => nios2_qsys_instruction_master_read,                            --                                       .read
			nios2_qsys_instruction_master_readdata       => nios2_qsys_instruction_master_readdata,                        --                                       .readdata
			nios2_qsys_instruction_master_readdatavalid  => nios2_qsys_instruction_master_readdatavalid,                   --                                       .readdatavalid
			jtag_uart_avalon_jtag_slave_address          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,         --            jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write            => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,           --                                       .write
			jtag_uart_avalon_jtag_slave_read             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,            --                                       .read
			jtag_uart_avalon_jtag_slave_readdata         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                                       .readdata
			jtag_uart_avalon_jtag_slave_writedata        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                                       .writedata
			jtag_uart_avalon_jtag_slave_waitrequest      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                                       .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      --                                       .chipselect
			mm_clock_crossing_bridge_0_s0_address        => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address,       --          mm_clock_crossing_bridge_0_s0.address
			mm_clock_crossing_bridge_0_s0_write          => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write,         --                                       .write
			mm_clock_crossing_bridge_0_s0_read           => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read,          --                                       .read
			mm_clock_crossing_bridge_0_s0_readdata       => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata,      --                                       .readdata
			mm_clock_crossing_bridge_0_s0_writedata      => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata,     --                                       .writedata
			mm_clock_crossing_bridge_0_s0_burstcount     => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount,    --                                       .burstcount
			mm_clock_crossing_bridge_0_s0_byteenable     => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable,    --                                       .byteenable
			mm_clock_crossing_bridge_0_s0_readdatavalid  => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid, --                                       .readdatavalid
			mm_clock_crossing_bridge_0_s0_waitrequest    => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest,   --                                       .waitrequest
			mm_clock_crossing_bridge_0_s0_debugaccess    => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess,   --                                       .debugaccess
			nios2_qsys_debug_mem_slave_address           => mm_interconnect_0_nios2_qsys_debug_mem_slave_address,          --             nios2_qsys_debug_mem_slave.address
			nios2_qsys_debug_mem_slave_write             => mm_interconnect_0_nios2_qsys_debug_mem_slave_write,            --                                       .write
			nios2_qsys_debug_mem_slave_read              => mm_interconnect_0_nios2_qsys_debug_mem_slave_read,             --                                       .read
			nios2_qsys_debug_mem_slave_readdata          => mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata,         --                                       .readdata
			nios2_qsys_debug_mem_slave_writedata         => mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata,        --                                       .writedata
			nios2_qsys_debug_mem_slave_byteenable        => mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable,       --                                       .byteenable
			nios2_qsys_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest,      --                                       .waitrequest
			nios2_qsys_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess,      --                                       .debugaccess
			onchip_mem_s1_address                        => mm_interconnect_0_onchip_mem_s1_address,                       --                          onchip_mem_s1.address
			onchip_mem_s1_write                          => mm_interconnect_0_onchip_mem_s1_write,                         --                                       .write
			onchip_mem_s1_readdata                       => mm_interconnect_0_onchip_mem_s1_readdata,                      --                                       .readdata
			onchip_mem_s1_writedata                      => mm_interconnect_0_onchip_mem_s1_writedata,                     --                                       .writedata
			onchip_mem_s1_byteenable                     => mm_interconnect_0_onchip_mem_s1_byteenable,                    --                                       .byteenable
			onchip_mem_s1_chipselect                     => mm_interconnect_0_onchip_mem_s1_chipselect,                    --                                       .chipselect
			onchip_mem_s1_clken                          => mm_interconnect_0_onchip_mem_s1_clken,                         --                                       .clken
			sdram_s1_address                             => mm_interconnect_0_sdram_s1_address,                            --                               sdram_s1.address
			sdram_s1_write                               => mm_interconnect_0_sdram_s1_write,                              --                                       .write
			sdram_s1_read                                => mm_interconnect_0_sdram_s1_read,                               --                                       .read
			sdram_s1_readdata                            => mm_interconnect_0_sdram_s1_readdata,                           --                                       .readdata
			sdram_s1_writedata                           => mm_interconnect_0_sdram_s1_writedata,                          --                                       .writedata
			sdram_s1_byteenable                          => mm_interconnect_0_sdram_s1_byteenable,                         --                                       .byteenable
			sdram_s1_readdatavalid                       => mm_interconnect_0_sdram_s1_readdatavalid,                      --                                       .readdatavalid
			sdram_s1_waitrequest                         => mm_interconnect_0_sdram_s1_waitrequest,                        --                                       .waitrequest
			sdram_s1_chipselect                          => mm_interconnect_0_sdram_s1_chipselect                          --                                       .chipselect
		);

	mm_interconnect_1 : component DE0_CV_QSYS_mm_interconnect_1
		port map (
			pll_outclk2_clk                                                 => pll_outclk2_clk,                                     --                                               pll_outclk2.clk
			mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                  -- mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset.reset
			transmitter_reset_n_reset_bridge_in_reset_reset                 => rst_controller_001_reset_out_reset,                  --                 transmitter_reset_n_reset_bridge_in_reset.reset
			mm_clock_crossing_bridge_0_m0_address                           => mm_clock_crossing_bridge_0_m0_address,               --                             mm_clock_crossing_bridge_0_m0.address
			mm_clock_crossing_bridge_0_m0_waitrequest                       => mm_clock_crossing_bridge_0_m0_waitrequest,           --                                                          .waitrequest
			mm_clock_crossing_bridge_0_m0_burstcount                        => mm_clock_crossing_bridge_0_m0_burstcount,            --                                                          .burstcount
			mm_clock_crossing_bridge_0_m0_byteenable                        => mm_clock_crossing_bridge_0_m0_byteenable,            --                                                          .byteenable
			mm_clock_crossing_bridge_0_m0_read                              => mm_clock_crossing_bridge_0_m0_read,                  --                                                          .read
			mm_clock_crossing_bridge_0_m0_readdata                          => mm_clock_crossing_bridge_0_m0_readdata,              --                                                          .readdata
			mm_clock_crossing_bridge_0_m0_readdatavalid                     => mm_clock_crossing_bridge_0_m0_readdatavalid,         --                                                          .readdatavalid
			mm_clock_crossing_bridge_0_m0_write                             => mm_clock_crossing_bridge_0_m0_write,                 --                                                          .write
			mm_clock_crossing_bridge_0_m0_writedata                         => mm_clock_crossing_bridge_0_m0_writedata,             --                                                          .writedata
			mm_clock_crossing_bridge_0_m0_debugaccess                       => mm_clock_crossing_bridge_0_m0_debugaccess,           --                                                          .debugaccess
			keys_s1_address                                                 => mm_interconnect_1_keys_s1_address,                   --                                                   keys_s1.address
			keys_s1_write                                                   => mm_interconnect_1_keys_s1_write,                     --                                                          .write
			keys_s1_readdata                                                => mm_interconnect_1_keys_s1_readdata,                  --                                                          .readdata
			keys_s1_writedata                                               => mm_interconnect_1_keys_s1_writedata,                 --                                                          .writedata
			keys_s1_chipselect                                              => mm_interconnect_1_keys_s1_chipselect,                --                                                          .chipselect
			leds_s1_address                                                 => mm_interconnect_1_leds_s1_address,                   --                                                   leds_s1.address
			leds_s1_write                                                   => mm_interconnect_1_leds_s1_write,                     --                                                          .write
			leds_s1_readdata                                                => mm_interconnect_1_leds_s1_readdata,                  --                                                          .readdata
			leds_s1_writedata                                               => mm_interconnect_1_leds_s1_writedata,                 --                                                          .writedata
			leds_s1_chipselect                                              => mm_interconnect_1_leds_s1_chipselect,                --                                                          .chipselect
			seg7_digits_s1_address                                          => mm_interconnect_1_seg7_digits_s1_address,            --                                            seg7_digits_s1.address
			seg7_digits_s1_write                                            => mm_interconnect_1_seg7_digits_s1_write,              --                                                          .write
			seg7_digits_s1_readdata                                         => mm_interconnect_1_seg7_digits_s1_readdata,           --                                                          .readdata
			seg7_digits_s1_writedata                                        => mm_interconnect_1_seg7_digits_s1_writedata,          --                                                          .writedata
			seg7_digits_s1_chipselect                                       => mm_interconnect_1_seg7_digits_s1_chipselect,         --                                                          .chipselect
			switches_s1_address                                             => mm_interconnect_1_switches_s1_address,               --                                               switches_s1.address
			switches_s1_readdata                                            => mm_interconnect_1_switches_s1_readdata,              --                                                          .readdata
			sysid_qsys_control_slave_address                                => mm_interconnect_1_sysid_qsys_control_slave_address,  --                                  sysid_qsys_control_slave.address
			sysid_qsys_control_slave_readdata                               => mm_interconnect_1_sysid_qsys_control_slave_readdata, --                                                          .readdata
			timer_s1_address                                                => mm_interconnect_1_timer_s1_address,                  --                                                  timer_s1.address
			timer_s1_write                                                  => mm_interconnect_1_timer_s1_write,                    --                                                          .write
			timer_s1_readdata                                               => mm_interconnect_1_timer_s1_readdata,                 --                                                          .readdata
			timer_s1_writedata                                              => mm_interconnect_1_timer_s1_writedata,                --                                                          .writedata
			timer_s1_chipselect                                             => mm_interconnect_1_timer_s1_chipselect,               --                                                          .chipselect
			transmitter_avalon_eln_address                                  => mm_interconnect_1_transmitter_avalon_eln_address,    --                                    transmitter_avalon_eln.address
			transmitter_avalon_eln_write                                    => mm_interconnect_1_transmitter_avalon_eln_write,      --                                                          .write
			transmitter_avalon_eln_read                                     => mm_interconnect_1_transmitter_avalon_eln_read,       --                                                          .read
			transmitter_avalon_eln_readdata                                 => mm_interconnect_1_transmitter_avalon_eln_readdata,   --                                                          .readdata
			transmitter_avalon_eln_writedata                                => mm_interconnect_1_transmitter_avalon_eln_writedata   --                                                          .writedata
		);

	irq_mapper : component DE0_CV_QSYS_irq_mapper
		port map (
			clk           => pll_outclk0_clk,                --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => nios2_qsys_irq_irq              --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_outclk2_clk,                    --       receiver_clk.clk
			sender_clk     => pll_outclk0_clk,                    --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_reset_out_reset,     --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_inv,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	irq_synchronizer_001 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_outclk2_clk,                    --       receiver_clk.clk
			sender_clk     => pll_outclk0_clk,                    --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_reset_out_reset,     --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_001_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver1_irq            --             sender.irq
		);

	irq_synchronizer_002 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_outclk2_clk,                    --       receiver_clk.clk
			sender_clk     => pll_outclk0_clk,                    --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_reset_out_reset,     --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_002_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver3_irq            --             sender.irq
		);

	rst_controller : component de0_cv_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,              -- reset_in0.reset
			reset_in1      => nios2_qsys_debug_reset_request_reset, -- reset_in1.reset
			clk            => pll_outclk0_clk,                      --       clk.clk
			reset_out      => rst_controller_reset_out_reset,       -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,   --          .reset_req
			reset_req_in0  => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	rst_controller_001 : component de0_cv_qsys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,              -- reset_in0.reset
			reset_in1      => nios2_qsys_debug_reset_request_reset, -- reset_in1.reset
			clk            => pll_outclk2_clk,                      --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,   -- reset_out.reset
			reset_req      => open,                                 -- (terminated)
			reset_req_in0  => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	rst_controller_002 : component de0_cv_qsys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,              -- reset_in0.reset
			reset_in1      => nios2_qsys_debug_reset_request_reset, -- reset_in1.reset
			clk            => open,                                 --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,   -- reset_out.reset
			reset_req      => open,                                 -- (terminated)
			reset_req_in0  => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_1_timer_s1_write_ports_inv <= not mm_interconnect_1_timer_s1_write;

	mm_interconnect_1_keys_s1_write_ports_inv <= not mm_interconnect_1_keys_s1_write;

	mm_interconnect_1_leds_s1_write_ports_inv <= not mm_interconnect_1_leds_s1_write;

	mm_interconnect_1_seg7_digits_s1_write_ports_inv <= not mm_interconnect_1_seg7_digits_s1_write;

	irq_synchronizer_receiver_inv(0) <= not transmitter_irq_eln_n_irq;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of DE0_CV_QSYS
